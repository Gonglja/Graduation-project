//module temp_tp();
//
//
//temp Temp(clk,nRST,Data,data1);
//
//endmodule
